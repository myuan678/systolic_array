


module pe_os #(
    localparam integer unsigned DIN_WIDTH = 8  ,
    localparam integer unsigned ACC_WIDTH = 32
)(
    input                       clk         ,
    input                       rst_n       ,
    input [DIN_WIDTH-1:0]       din_row     ,
    input [DIN_WIDTH-1:0]       din_col     ,

);
    
endmodule